* C:\Users\saisr\eSim-Workspace\parity_gen\parity_gen.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 5/14/2021 8:17:52 AM

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
U2  Net-_U2-Pad1_ Net-_U2-Pad2_ Net-_U2-Pad3_ Net-_U2-Pad4_ Net-_U2-Pad5_ parity_gen		
U6  in1 in2 in3 in4 Net-_U2-Pad1_ Net-_U2-Pad2_ Net-_U2-Pad3_ Net-_U2-Pad4_ adc_bridge_4		
U7  Net-_U2-Pad5_ out dac_bridge_1		
v1  in1 GND pulse		
v2  in2 GND pulse		
v3  in3 GND pulse		
v4  in4 GND pulse		
R1  out GND resistor		
U5  in1 plot_v1		
U4  in2 plot_v1		
U3  in3 plot_v1		
U1  in4 plot_v1		
U8  out plot_v1		

.end
